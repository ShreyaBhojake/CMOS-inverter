magic
tech sky130A
timestamp 1725783045
<< nwell >>
rect -250 400 50 890
<< nmos >>
rect -105 250 -90 350
<< pmos >>
rect -105 445 -90 655
<< ndiff >>
rect -150 340 -105 350
rect -150 260 -140 340
rect -120 260 -105 340
rect -150 250 -105 260
rect -90 340 -45 350
rect -90 260 -75 340
rect -55 260 -45 340
rect -90 250 -45 260
<< pdiff >>
rect -205 645 -105 655
rect -205 455 -195 645
rect -125 455 -105 645
rect -205 445 -105 455
rect -90 645 10 655
rect -90 455 -70 645
rect 0 455 10 645
rect -90 445 10 455
<< ndiffc >>
rect -140 260 -120 340
rect -75 260 -55 340
<< pdiffc >>
rect -195 455 -125 645
rect -70 455 0 645
<< psubdiff >>
rect -165 205 -25 220
rect -165 165 -150 205
rect -40 165 -25 205
rect -165 150 -25 165
<< nsubdiff >>
rect -225 835 25 845
rect -225 830 -145 835
rect -120 830 25 835
rect -225 770 -200 830
rect 0 770 25 830
rect -225 760 -145 770
rect -120 760 25 770
rect -225 755 25 760
<< psubdiffcont >>
rect -150 165 -40 205
<< nsubdiffcont >>
rect -145 830 -120 835
rect -200 770 0 830
rect -145 760 -120 770
<< poly >>
rect -105 655 -90 720
rect -105 425 -90 445
rect -180 415 -90 425
rect -180 390 -165 415
rect -140 390 -90 415
rect -180 380 -90 390
rect -65 415 -10 425
rect -65 390 -50 415
rect -25 390 -10 415
rect -65 380 -10 390
rect -105 350 -90 380
rect -105 235 -90 250
<< polycont >>
rect -165 390 -140 415
rect -50 390 -25 415
<< locali >>
rect -225 835 25 845
rect -225 830 -145 835
rect -70 830 25 835
rect -225 770 -200 830
rect 0 770 25 830
rect -225 760 -145 770
rect -70 760 25 770
rect -225 755 25 760
rect -200 655 -130 755
rect -205 645 -110 655
rect -205 455 -195 645
rect -125 455 -110 645
rect -205 445 -110 455
rect -85 645 10 655
rect -85 455 -70 645
rect 0 455 10 645
rect -85 445 10 455
rect -85 425 -45 445
rect -180 415 -125 425
rect -180 390 -165 415
rect -140 390 -125 415
rect -180 380 -125 390
rect -85 415 -10 425
rect -85 390 -50 415
rect -25 390 -10 415
rect -85 380 -10 390
rect -150 340 -110 350
rect -150 260 -140 340
rect -120 260 -110 340
rect -150 250 -110 260
rect -85 340 -45 380
rect -85 260 -75 340
rect -55 260 -45 340
rect -85 250 -45 260
rect -145 225 -110 250
rect -145 215 -120 225
rect -160 205 -120 215
rect -65 205 -30 215
rect -160 165 -150 205
rect -40 165 -30 205
rect -160 155 -120 165
rect -145 150 -120 155
rect -65 155 -30 165
<< viali >>
rect -145 830 -120 835
rect -120 830 -70 835
rect -145 770 -70 830
rect -145 760 -120 770
rect -120 760 -70 770
rect -165 390 -140 415
rect -50 390 -25 415
rect -120 205 -65 225
rect -120 165 -65 205
rect -120 150 -65 165
<< metal1 >>
rect -360 835 165 845
rect -360 760 -145 835
rect -70 760 165 835
rect -360 755 165 760
rect -360 415 -125 425
rect -360 390 -165 415
rect -140 390 -125 415
rect -360 380 -125 390
rect -85 415 185 425
rect -85 390 -50 415
rect -25 390 185 415
rect -85 380 185 390
rect -335 225 190 235
rect -335 150 -120 225
rect -65 150 190 225
rect -335 145 190 150
<< labels >>
rlabel metal1 105 800 105 800 1 vdd
rlabel metal1 105 185 105 185 1 vss
rlabel metal1 160 390 175 415 1 out
rlabel metal1 -350 390 -335 415 1 in
<< end >>
