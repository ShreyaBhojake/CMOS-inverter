magic
tech sky130A
timestamp 1725780265
<< nwell >>
rect -250 400 50 890
<< nmos >>
rect -105 250 -90 350
<< pmos >>
rect -105 445 -90 655
<< ndiff >>
rect -150 340 -105 350
rect -150 260 -140 340
rect -120 260 -105 340
rect -150 250 -105 260
rect -90 340 -45 350
rect -90 260 -75 340
rect -55 260 -45 340
rect -90 250 -45 260
<< pdiff >>
rect -205 645 -105 655
rect -205 455 -195 645
rect -125 455 -105 645
rect -205 445 -105 455
rect -90 645 10 655
rect -90 455 -70 645
rect 0 455 10 645
rect -90 445 10 455
<< ndiffc >>
rect -140 260 -120 340
rect -75 260 -55 340
<< pdiffc >>
rect -195 455 -125 645
rect -70 455 0 645
<< psubdiff >>
rect -165 205 -25 220
rect -165 165 -150 205
rect -40 165 -25 205
rect -165 150 -25 165
<< nsubdiff >>
rect -225 830 25 845
rect -225 770 -200 830
rect 0 770 25 830
rect -225 755 25 770
<< psubdiffcont >>
rect -150 165 -40 205
<< nsubdiffcont >>
rect -200 770 0 830
<< poly >>
rect -105 655 -90 720
rect -105 350 -90 445
rect -105 235 -90 250
<< locali >>
rect -225 830 25 845
rect -225 770 -200 830
rect 0 770 25 830
rect -225 755 25 770
rect -205 645 -110 655
rect -205 455 -195 645
rect -125 455 -110 645
rect -205 445 -110 455
rect -85 645 10 655
rect -85 455 -70 645
rect 0 455 10 645
rect -85 445 10 455
rect -150 340 -110 350
rect -150 260 -140 340
rect -120 260 -110 340
rect -150 250 -110 260
rect -85 340 -45 350
rect -85 260 -75 340
rect -55 260 -45 340
rect -85 250 -45 260
rect -160 205 -30 215
rect -160 165 -150 205
rect -40 165 -30 205
rect -160 155 -30 165
<< end >>
